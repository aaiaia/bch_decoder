`ifndef M_SBS_HARD_T3_COMB_PIPELINED
`define M_SBS_HARD_T3_COMB_PIPELINED

`include "00_GF_mult/gf_10/comb/GF_Mult_2_10_comb.v"

module mSBS_t3_comb_pipelined
(
    clk,
    in_ctr_Srst,
    in_ctr_en,

    synd1,
    synd3,
    synd5,

    out_deg2_A,
    out_deg2_B,
//    out_deg2_C,
    //out_deg2_R,

    out_deg3_A,
    out_deg3_B,
    out_deg3_C,
    out_deg3_R
);
    parameter   OUTTER_NAME = "";
    parameter   MODULE_NAME = "mSBS_t3_comb";
        localparam  DESIGN_NAME = "mSBS_t3_comb";

    parameter           GF_LEN  =   10;

    parameter   SYN_TEST    =   0;
    
    initial begin
        $display("!!! in) %s !!!", OUTTER_NAME);
        $display("!!! %s !!!", MODULE_NAME);
        $display("!!! %s !!!", DESIGN_NAME);

        $display("GF_LEN=%d", GF_LEN);
        $display("SYN_TEST=%d", SYN_TEST);
    end

    input                       clk;

    input                       in_ctr_Srst;
    input                       in_ctr_en;


    input       [GF_LEN-1:0]    synd1;
    input       [GF_LEN-1:0]    synd3;
    input       [GF_LEN-1:0]    synd5;

    output      [GF_LEN-1:0]    out_deg2_A;
    output      [GF_LEN-1:0]    out_deg2_B;
//    output      [GF_LEN-1:0]    out_deg2_C;
    //output      [GF_LEN-1:0]    out_deg2_R;

    output      [GF_LEN-1:0]    out_deg3_A;
    output      [GF_LEN-1:0]    out_deg3_B;
    output      [GF_LEN-1:0]    out_deg3_C;
    output      [GF_LEN-1:0]    out_deg3_R;


    wire        [GF_LEN-1:0]    synd1p2;
    wire        [GF_LEN-1:0]    synd1p3;

    wire        [GF_LEN-1:0]    synd1p2_synd3;

    wire        [GF_LEN-1:0]    Cp2;
    wire        [GF_LEN-1:0]    synd1_A;

    wire        [GF_LEN-1:0]    t2_R;
    wire        [GF_LEN-1:0]    t2_A;
    wire        [GF_LEN-1:0]    t2_B;
//    wire        [GF_LEN-1:0]    t2_C;

    wire        [GF_LEN-1:0]    t3_R;
    wire        [GF_LEN-1:0]    t3_A;
    wire        [GF_LEN-1:0]    t3_B;
    wire        [GF_LEN-1:0]    t3_C;


    reg         [GF_LEN-1:0]    pipe_s1p2s3_s5;
    reg         [GF_LEN-1:0]    pipe_s1p2;
    reg         [GF_LEN-1:0]    pipe_s1p3_s3;
    reg         [GF_LEN-1:0]    pipe_s1;

    always@(posedge clk) begin
        if(in_ctr_Srst) pipe_s1 <= {(GF_LEN){1'b0}};
        else if(in_ctr_en) pipe_s1 <= synd1;
        else pipe_s1 <= pipe_s1;
    end



    /* if error less than 3 start */
    assign t2_R = pipe_s1p3_s3;
    always@(posedge clk) begin
        if(in_ctr_Srst)pipe_s1p3_s3 <= {(GF_LEN){1'b0}};
        else if(in_ctr_en) pipe_s1p3_s3 <= t3_C;
        else pipe_s1p3_s3 <= pipe_s1p3_s3; 
    end
    assign t2_A = synd1p2;
    assign t2_B = pipe_s1;
    //assign t2_C = 0;
    /* if error less than 3 end */

    /* base start */
    GF_Mult_2_10_comb synd1_pow_2
    (
        .out(synd1p2),
        .a(synd1),
        .b(synd1)
    );

    GF_Mult_2_10_comb synd1_pow_3
    (
        .out(synd1p3),
        .a(synd1p2),
        .b(synd1)
    );
    /* base end */


    /* coeffi t3 A start */
    GF_Mult_2_10_comb mul_synd1p2_synd3
    (
        .out(synd1p2_synd3),
        .a(synd1p2),
        .b(synd3)
    );

    always@(posedge clk) begin
        if(in_ctr_Srst) pipe_s1p2s3_s5 <= {(GF_LEN){1'b0}};
        else if(in_ctr_en)  pipe_s1p2s3_s5 <= t3_A;
        else            pipe_s1p2s3_s5 <= pipe_s1p2s3_s5;
    end
    assign t3_A = synd1p2_synd3 ^ synd5;
    /* coeffi t3 A end */


    /* coeffi t3 C start */
    assign t3_C = synd1p3 ^ synd3;
    /* coeffi t3 C end */


    /* coeffi t3 B start */
    GF_Mult_2_10_comb mul_C_synd1
    (
        .out(t3_B),
        .a(pipe_s1p3_s3),
        .b(pipe_s1)
    );
    /* coeffi t3 B end */


    /* coeffi t3 R start */
    /* coeffi t3 R1*/
    GF_Mult_2_10_comb mul_C_pow2
    (
        .out(Cp2),
        .a(pipe_s1p3_s3),
        .b(pipe_s1p3_s3)
    );

    /* coeffi t3 R2 */
    GF_Mult_2_10_comb mul_synd1_A
    (
        .out(synd1_A),
        .a(pipe_s1p2s3_s5),
        .b(pipe_s1)
    );

    assign t3_R = Cp2 ^ synd1_A;
    /* coeffi t3 R end */
  
    /* error less than 3 detector */
    //assign detector = |pipe_s1p3_s3;

    //assign R = detector ? t3_R : t2_R;
    //assign A = detector ? pipe_s1p2s3_s5 : t2_A;
    //assign B = detector ? t3_B : t2_B;
    //assign C = detector ? pipe_s1p3_s3 : t2_C;

    generate
        if(!SYN_TEST) begin : gen_not_syn_test
            //assign  out_deg2_R = t2_R;
            always@(posedge clk) begin
                if(in_ctr_Srst)     pipe_s1p2 <= {(GF_LEN){1'b0}};
                else if(in_ctr_en)  pipe_s1p2 <= t2_A;
                else                pipe_s1p2 <= pipe_s1p2;
            end
            //assign  out_deg2_A = t2_A;
            assign  out_deg2_A = pipe_s1p2;
            assign  out_deg2_B = t2_B;
//            assign  out_deg2_C = t2_C;
                      
            assign  out_deg3_R = t3_R;
            assign  out_deg3_A = pipe_s1p2s3_s5;
            assign  out_deg3_B = t3_B;
            assign  out_deg3_C = pipe_s1p3_s3;
        end
        else begin
            reg [GF_LEN - 1 : 0]    buf_deg3_R;
            reg [GF_LEN - 1 : 0]    buf_deg3_A;
            reg [GF_LEN - 1 : 0]    buf_deg3_B;
            reg [GF_LEN - 1 : 0]    buf_deg3_C;

            reg [GF_LEN - 1 : 0]    buf_deg2_R;
            reg [GF_LEN - 1 : 0]    buf_deg2_A;
            reg [GF_LEN - 1 : 0]    buf_deg2_B;
            reg [GF_LEN - 1 : 0]    buf_deg2_C;
                                              
            always@(posedge clk) begin
                buf_deg3_R <= t2_R;
                buf_deg3_A <= t2_A;
                buf_deg3_B <= t2_B;
//                buf_deg3_C <= t2_C;
                                 
                buf_deg2_R <= t3_R; 
                buf_deg2_A <= pipe_s1p2s3_s5;
                buf_deg2_B <= t3_B;
                buf_deg2_C <= pipe_s1p3_s3;
            end    


            //assign  out_deg2_R = buf_deg2_R;
            assign  out_deg2_A = buf_deg2_A;
            assign  out_deg2_B = buf_deg2_B;
//            assign  out_deg2_C = buf_deg2_C;
                                   
            assign  out_deg3_R = buf_deg3_R;
            assign  out_deg3_A = buf_deg3_A;
            assign  out_deg3_B = buf_deg3_B;
            assign  out_deg3_C = buf_deg3_C;


        end
    endgenerate







endmodule

`endif
